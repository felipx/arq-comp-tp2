//! @title TRANSMITTER
//! @file transmitter.v
//! @author Felipe Montero Bruni
//! @date 10-2023
//! @version 0.1

module transmitter #(
    parameters
) (
    ports
);
    
endmodule